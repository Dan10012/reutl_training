//////////////////////////////////////////////////////////////////
///
/// Project Name: 	avalon_enforced
///
/// File Name: 		avalon_enforced_pack.sv
///
//////////////////////////////////////////////////////////////////
///
/// Author: 		Reut Lev
///
/// Date Created: 	26.3.2020
///
/// Company: 		----
///
//////////////////////////////////////////////////////////////////
///
/// Description: 	?????
///
//////////////////////////////////////////////////////////////////

package avalon_enforced_pack;
	
	typedef enum {
		WAIT_FOR_MESSAGE,
		RECIEVE_MASSAGE
	} avalon_enforced_sm_t;

endpackage